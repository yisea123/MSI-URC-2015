-- https://www.eewiki.net/display/LOGIC/Serial+Peripheral+Interface+%28SPI%29+Slave+%28VHDL%29